module RAM(
    input logic[31:0] address,
    input logic clk,
    output logic[31:0] read_data,
    input logic[31:0] write_data,
    input logic write_enable
);

reg[31:0] memory [4999:0];
integer i;
initial begin
    for(i = 0; i < 5000; i++) memory[i] = 0;

    $readmemb("test1.txt", memory);
    for (i = 0; i < 24; i++) begin
        $display("%h: %h", (i*4), memory[i]);
    end


end

always_ff @(posedge clk)begin
    if(write_enable) memory[address/4] <= write_data;
    read_data <= memory[address/4];
end

endmodule